//***************************************
// Parameter definitions
//***************************************

parameter ROWS=16;	//Quantity of rows in memory array
parameter COLS=16;	//Quantity of columns in memory array
