parameter ROWS=2;
parameter COLS=8;
