//***************************************
// Parameter definitions
//***************************************

parameter ROWS=8;	//Quantity of rows in memory array
parameter COLS=8;	//Quantity of columns in memory array
