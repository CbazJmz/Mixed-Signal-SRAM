module nmospass
(
	inout wire d,
	inout wire s,
	input wire g
);

	nmos(d,s,g);

	endmodule
