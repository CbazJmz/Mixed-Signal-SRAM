parameter ROWS=8;
parameter COLS=8;
